module UATransmit(
  input   Clock,
  input   Reset,

  input   [7:0] DataIn,
  input         DataInValid,
  output        DataInReady,

  output        SOut
);
    // for log2 function
    `include "util.vh"

    //--|Parameters|--------------------------------------------------------------
    parameter   ClockFreq         =   100_000_000;
    parameter   BaudRate          =   115_200;

    // See diagram in the lab guide
    localparam  SymbolEdgeTime    =   ClockFreq / BaudRate;
    localparam  ClockCounterWidth =   log2(SymbolEdgeTime);

    // Copy your UART transmitter implementation from Lab 6 to here.

endmodule
