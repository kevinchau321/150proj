/**
 * Top-level module for the RISCV processor.
 * This should contain instantiations of your datapath and control unit.
 * For CP1, the imem and dmem should be instantiated in this top-level module.
 * For CP2 and CP3, the memories are moved to a different module (Memory150),
 * and connected to the datapath via memory ports in the RISC I/O interface.
 *
 * CS150 Fall 14. Template written by Simon Scott.
 */
module Riscv150(
    input clk,
    input rst,
    input stall,

    // Ports for UART that go off-chip to UART level shifter
    input FPGA_SERIAL_RX,
    output FPGA_SERIAL_TX

    // Memory system ports
    // Only used for checkpoint 2 and 3
`ifdef CS150_CHKPNT_2_OR_3
    ,
    output [31:0] dcache_addr,
    output [31:0] icache_addr,
    output [3:0] dcache_we,
    output [3:0] icache_we,
    output dcache_re,
    output icache_re,
    output [31:0] dcache_din,
    output [31:0] icache_din,
    input [31:0] dcache_dout,
    input [31:0] instruction
`endif

    // Graphics ports
    // Only used for checkpoint 3
`ifdef CS150_CHKPNT_3
    ,
    output [31:0]  bypass_addr,
    output [31:0]  bypass_din,
    output [3:0]   bypass_we,

    input          filler_ready,
    input          line_ready,
    output  [23:0] filler_color,
    output         filler_valid,
    output  [31:0] line_color,
    output  [9:0]  line_point,
    output         line_color_valid,
    output         line_x0_valid,
    output         line_y0_valid,
    output         line_x1_valid,
    output         line_y1_valid,
    output         line_trigger
`endif
);


    wire [7:0] UARTtoWB;
    // Instantiate the instruction memory here (checkpoint 1 only)
    imem_blk_ram(.clka(clk),
		.ena(),
		.wea(),
		.addra(),
		.dina(),
		.clkb(),
		.addrb(),
		.doutb());

    // Instantiate the data memory here (checkpoint 1 only)
    dmem_blk_ram(.clka(clk), 
		.ena(),
		.wea(),
		.addra(),
		.dina(),
		.douta());
    // Instantiate your control unit here
   //ControlUnit control(
//		.UART_out(UARTtoWB)
//);
    // Instantiate your datapath here
   Datapath datapath ();
   UART uart(
	.SIn(FPGA_SERIAL_RX),
	.SOut(FPGA_SERIAL_TX),	
	.DataOut(UARTtoWB));
   
   
endmodule
