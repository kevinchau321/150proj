module asmtest(input clk, input rst, input [29:0] addr, output reg [31:0] inst);
reg [29:0] addr_r;
always @(posedge clk)
begin
addr_r <= (rst) ? (30'b0) : (addr);
end
always @(*)
begin
case(addr_r)
30'h00000000: inst = 32'h93030000;
30'h00000001: inst = 32'hb7000010;
30'h00000002: inst = 32'h93800002;
30'h00000003: inst = 32'h37b1ad1e;
30'h00000004: inst = 32'h1301f10e;
30'h00000005: inst = 32'h37050010;
30'h00000006: inst = 32'h23201500;
30'h00000007: inst = 32'h23222500;
30'h00000008: inst = 32'h83250500;
30'h00000009: inst = 32'h03264500;
30'h0000000a: inst = 32'h6398b000;
30'h0000000b: inst = 32'h93831300;
30'h0000000c: inst = 32'h6314c100;
30'h0000000d: inst = 32'h6f008004;
30'h0000000e: inst = 32'h13026004;
30'h0000000f: inst = 32'hef000007;
30'h00000010: inst = 32'h13021006;
30'h00000011: inst = 32'hef008006;
30'h00000012: inst = 32'h13029006;
30'h00000013: inst = 32'hef000006;
30'h00000014: inst = 32'h1302c006;
30'h00000015: inst = 32'hef008005;
30'h00000016: inst = 32'h1302a003;
30'h00000017: inst = 32'hef000005;
30'h00000018: inst = 32'h13020002;
30'h00000019: inst = 32'hef008004;
30'h0000001a: inst = 32'h13820303;
30'h0000001b: inst = 32'hef000004;
30'h0000001c: inst = 32'h1302a000;
30'h0000001d: inst = 32'hef008003;
30'h0000001e: inst = 32'h6f000003;
30'h0000001f: inst = 32'h13020005;
30'h00000020: inst = 32'hef00c002;
30'h00000021: inst = 32'h13021006;
30'h00000022: inst = 32'hef004002;
30'h00000023: inst = 32'h13023007;
30'h00000024: inst = 32'hef00c001;
30'h00000025: inst = 32'h13023007;
30'h00000026: inst = 32'hef004001;
30'h00000027: inst = 32'h1302a000;
30'h00000028: inst = 32'hef00c000;
30'h00000029: inst = 32'h6f004000;
30'h0000002a: inst = 32'h6f000000;
30'h0000002b: inst = 32'h37010080;
30'h0000002c: inst = 32'h83210100;
30'h0000002d: inst = 32'h93f11100;
30'h0000002e: inst = 32'he38a01fe;
30'h0000002f: inst = 32'h23244100;
30'h00000030: inst = 32'h67800000;
default:      inst = 32'h00000000;
endcase
end
endmodule
